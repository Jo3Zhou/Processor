library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity dual_port_mem is --memory for storing and reading instruction & data
    Port ( clk : in STD_LOGIC;
           wen : in STD_LOGIC;
           ins_add : in STD_LOGIC_VECTOR (6 downto 0);
           ins : out STD_LOGIC_VECTOR (31 downto 0);
           data_add : in STD_LOGIC_VECTOR (6 downto 0);
           data_in : in STD_LOGIC_VECTOR (31 downto 0);
           data_out : out STD_LOGIC_VECTOR (31 downto 0));
end dual_port_mem;

architecture Behavioral of dual_port_mem is

type ram_array is array (0 to 127) of STD_LOGIC_VECTOR(31 downto 0);
    signal ram:ram_array:=(
    0  => B"00000000000000000000000000000000",  --instruction 0
    1  => B"10000100000001111100000000001111",
    2  => B"11000000000001111111110111100000",
    3  => B"00011000000000000111110000011111",
    4  => B"00010000000000000000000000000001",
    5  => B"00100000000000000000000000100001",
    6  => B"11001100000000000001011111100000",
    7  => B"10011000000000000000001111100001",
    8  => B"00100000000000000000000000100001",
    9  => B"00100100000000000000001111111111",
    10 => B"11011100000001111111000000000000",
    11 => B"10000100000000000100000000000010",
    12 => B"01010100000000000001000000011110",
    13 => B"10001000000000000000001111000011", 
    14 => B"10001100000000000000111111000100",
    15 => B"01011011111111111111110000011101",
    16 => B"10000000000000000000000000000111",
    17 => B"01010000000000000100001110100101",
    18 => B"01010000000000000000010010000110",
    19 => B"11000000000000000000100011000000",
    20 => B"00010000000000000001110001100111",
    21 => B"01100100000000000000010010000100",
    22 => B"01100000000000000000010001100011",
    23 => B"00100100000000000000000010100101",
    24 => B"11000100000001111110100010100000",
    25 => B"10010100000000000000000000000111",
    26 => B"01101000000000000010010011100111",
    27 => B"01101100000000000000110011100111",
    28 => B"01000000000000000000000011101000",
    29 => B"01001100000000000111010100001000",
    30 => B"00010100000000000010000011101001",
    31 => B"00011100000000000000010100101010",
    32 => B"11010000000000000010010101000000",
    33 => B"11011000000000000010000101000000",
    34 => B"00011000000000000000100101001011",
    35 => B"11010100000000000001100101100000",
    36 => B"01001000000000000001110101101100",
    37 => B"10011100000000000000010000001100",
    38 => B"01000100000000000011000101101100",
    39 => B"11001000000000000000110110000000",
    40 => B"11011100000000000000000000000000",
    41 => B"11011100000000000000000000000000",
    42 => B"10010100000001111110000000000111",
    43 => B"11011100000000000000000000000000",
    
    others => B"00000000000000000000000000000000");

begin    
    process (clk)   --Synchronous write
    begin
        if(rising_edge(clk))then
            if(wen = '1')then
            ram(to_integer(unsigned(data_add))) <= data_in;
            end if;
        end if;
    end process;
    
    ins <= ram(to_integer(unsigned(ins_add)));  --Asynchronous read
    
    data_out <= ram(to_integer(unsigned(data_add))); 

    
end Behavioral;
